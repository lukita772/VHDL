library ieee;
use ieee.std_logic_1164.all;

entity myGenCnt is
	port(
		clk: in std_logic;
		rst: in std_logic;
		q: out std_logic_vector(2 downto 0)
	);
end myGenCnt;

architecture arch_myGenCnt of myGenCnt is

begin

end arch_myGenCnt;
